Library ieee;
Use ieee.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY tb_Sign_Extension_Unit IS
GENERIC(N:INTEGER:=16;
M:INTEGER:=32);
END ENTITY;


ARCHITECTURE ARC OF tb_Sign_Extension_Unit IS
COMPONENT Sign_Extension_Unit IS
GENERIC(N:INTEGER:=16;
M:INTEGER:=32);
PORT(INPUT: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
OUTPUT: OUT STD_LOGIC_VECTOR(M-1 DOWNTO 0)
);
END COMPONENT;

SIGNAL tINPUT: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
SIGNAL tOUTPUT: STD_LOGIC_VECTOR(M-1 DOWNTO 0);

--clock signal and clock_period constant
SIGNAL tCLK: STD_LOGIC;
CONSTANT CLOCK_PERIOD: time:=100 ps;
--HERE COME COMPONENTS DECLARATIONS, SIGNALS,TYPES,CONSTANTS--
BEGIN
--PORT MAPPINGS COMES HERE
Sign_Extension_Unit_COMP: Sign_Extension_Unit PORT MAP(tINPUT,tOUTPUT);
PROCESS (TCLK)
BEGIN
--PROCESS CODE HERE
END PROCESS;

--The Clock Process: a process used for the testbench to not even have to enter this
tCLK<=NOT tCLK AFTER CLOCK_PERIOD/2;
--PORT MAP HERE--
PROCESS(Tclk)
BEGIN
tCLK<=NOT tCLK AFTER CLOCK_PERIOD/2;
END PROCESS;
--OTHER ARCHITECTURAL COMPONENTS

END ARC;
