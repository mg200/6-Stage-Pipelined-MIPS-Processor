Library ieee;
Use ieee.std_logic_1164.all;

ENTITY mux_4x1 IS
GENERIC(N:INTEGER:=16);
PORT(
I0,I1,I2,I3: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
Y:OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END ENTITY;

---STRUCTURAL DESIGN USING 2X1 MUXES
ARCHITECTURE ARC_BY_2X1_MUXES OF mux_4x1 IS
COMPONENT MUX_2X1_GENERIC IS
GENERIC(N: INTEGER:=16);
PORT(
I0,I1: IN STD_LOGIC_VECTOR( N-1 DOWNTO 0);
S: IN STD_LOGIC;
Y: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END COMPONENT;

SIGNAL tY0,tY1,tY2: STD_LOGIC_VECTOR(N-1 DOWNTO 0);

BEGIN
M0: MUX_2X1_GENERIC GENERIC MAP(N) PORT MAP(I0,I1,S(0),tY0);
M1: MUX_2X1_GENERIC GENERIC MAP(N) PORT MAP(I2,I3,S(0),tY1);
M2: MUX_2X1_GENERIC GENERIC MAP(N) PORT MAP(tY0,tY1,S(1),Y);
END ARC_BY_2X1_MUXES;
