Library ieee;
Use ieee.std_logic_1164.all;

ENTITY IntegratedUnit IS

PORT(

CLK: INOUT STD_LOGIC;--:='0';
EN: IN STD_LOGIC:='1';
RST: IN STD_LOGIC:='0'
-- output: out std_logic_vector(3 downto 0);
-- output2: out std_logic_vector(2 downto 0)
);

END IntegratedUnit;

ARCHITECTURE ARC OF IntegratedUnit IS




COMPONENT PC IS
GENERIC(N: INTEGER:=8);
PORT(CLK: IN STD_LOGIC:='1';
COUNT: inOUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
EN: IN STD_LOGIC:='1';
RST: IN STD_LOGIC:='0'
);
END COMPONENT;

COMPONENT RAM_GENERIC IS
GENERIC(
ADD_WIDTH: INTEGER:=8;
 DATA_WIDTH:INTEGER:=16);
PORT(
DATA_IN: IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
-- ADDRESS: IN STD_LOGIC_VECTOR(log2_unsigned(ADD_WIDTH)-1 DOWNTO 0);
ADDRESS: IN STD_LOGIC_VECTOR(ADD_WIDTH-1 DOWNTO 0);
READ_WRITE: IN STD_LOGIC:='1';--DEFAULT IS 1 TO WRITE
CLK: IN STD_LOGIC;
DATAOUT: OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
);
END COMPONENT;
COMPONENT A_REGISTER IS
GENERIC(N: INTEGER:=8);
PORT( 
D: IN STd_LOGIC_VECTOR(N-1 DOWNTO 0);
CLK,EN,RST: IN STD_LOGIC;
Q: OUT  STd_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;

COMPONENT CONTROLLER IS
PORT(
CLK: IN STD_LOGIC;
INPUT: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
ALU_OPERATION: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
CIN: OUT STD_LOGIC;
WRITE_EN: OUT STD_LOGIC
--READ_EN: OUT STD_LOGIC
);
END COMPONENT;


-- COMPONENT array_registerfile is
--     generic(N: INTEGER:=8);
--     PORT(
--         RESET : IN STD_LOGIC;
--         CLK: IN STd_LOGIC;
--         WRITE_ENABLE: IN STD_LOGIC;--_VECTOR(N-1 DOWNTO 0);
--         READ_ADD1, READ_ADD2: IN STd_LOGIC_VECTOR(2 DOWNTO 0);
--         WRITE_ADD: IN  STd_LOGIC_VECTOR(2 DOWNTO 0);
--         READ_PORT1, READ_PORT2: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
--         WRITE_PORT: IN STD_LOGIC_VECTOR (N-1 DOWNTO 0)
--         );
-- end COMPONENT;

COMPONENT array_registerfile is
    generic(N: INTEGER:=3);
    PORT(
        RESET : IN STD_LOGIC;
        CLK: IN STd_LOGIC;
WRITE_ENABLE: IN STD_LOGIC;--_VECTOR(N-1 DOWNTO 0);
        READ_ADD1, READ_ADD2: IN STd_LOGIC_VECTOR(N-1 DOWNTO 0);
        WRITE_ADD: IN  STd_LOGIC_VECTOR(N-1 DOWNTO 0);
        READ_PORT1, READ_PORT2: OUT STd_LOGIC_VECTOR((2**N)-1 DOWNTO 0);
        WRITE_PORT: IN STd_LOGIC_VECTOR ((2**N)-1 DOWNTO 0)
        );
end COMPONENT;


COMPONENT ALU IS
GENERIC(N:INTEGER:=8);
PORT(A,B: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
SELECTION: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
CIN: IN STD_LOGIC;
F: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
COUT: OUT STD_LOGIC
);

END COMPONENT;
--end of components
signal tclk: std_logic;
signal PC_ADD: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL T_INST,T_FETCH: STD_LOGIC_VECTOR(15 DOWNTO 0):=(others=>'0');
SIGNAL CONT_WRITE_EN: STD_LOGIC;
SIGNAL CONT_ALU_OP: STD_lOGIC_VECTOR(3 DOWNTO 0);
SIGNAL T_CIN: STD_LOGIC;
--REGISTER FILE SIGNALS 
SIGNAL tREADPORT1, tREADPORT2: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL tWRITE_PORT: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL tWRITEBACK_ADDRESS: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL DecExc_input: STD_LOGIC_VECTOR(24 DOWNTO 0);
---WRITE
SIGNAL WRITEBACK_ENABLE: STD_LOGIC;

--ALU SIGNALS
SIGNAL t_FETCH_EXECUTE: STD_LOGIC_VECTOR(24 DOWNTO 0);
SIGNAL tALU_OUTPUT: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL tALU_COUT: STD_LOGIC;

--WRITEBACK REGISTER
SIGNAL tWRITE_BACK_REGISTER: STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL WriteBack_Input: STD_LOGIC_VECTOR(11 DOWNTO 0);



-- CONSTANT CLOCK_PERIOD:TIME:= 100 ns;
BEGIN
-- CLK<=NOT CLK AFTER CLOCK_PERIOD/2;

--PC PORT MAP
PC_component: pc port map(CLK,PC_ADD,EN,RST);
--INSTRUCTION CACHE MEMORY PORT MAP--NOTE IT IS READ-ONLY SO WRITING IS DISENABLED
Inst_Cache_Component: ram_generic generic map(8,16) port map(X"0000",PC_ADD,'0',CLK,T_INST);
--Fetch_Decode Buffer PORT MAP
Fetch_Decode: A_REGISTER GENERIC MAP(16) PORT MAP(T_INST,clk,EN,rst,T_FETCH);
--CONTROLLER PORT MAP
CONT: CONTROLLER PORT MAP(CLK,T_FETCH(15 DOWNTO 13),CONT_ALU_OP,T_CIN,CONT_WRITE_EN);

--register file PORT MAP
register_file: ARRAY_REGISTERFILE PORT MAP(RST,CLK,WRITEBACK_ENABLE,T_FETCH(12 DOWNTO 10),
T_FETCH(9 DOWNTO 7),tWRITEBACK_ADDRESS,tREADPORT1,tREADPORT2,tWRITE_PORT);


--the output signal of the Fetch_Decode unit 
DecExc_input<=tREADPORT1&tREADPORT2&CONT_ALU_OP&T_FETCH(6 DOWNTO 4)&CONT_WRITE_EN&T_CIN;

--DECODE_EXECUTE_REGISTER PORT MAP
DECODE_EXECUTE_REGISTER: A_REGISTER GENERIC MAP(25) PORT MAP(DecExc_input,CLK,EN,RST,T_FETCH_EXECUTE);

--ALU PORT MAP
ALU_instance: ALU PORT MAP(T_fetch_execute(24 downto 17), t_fetch_execute(16 downto 9),
t_FETCH_EXECUTE(8 DOWNTO 5),T_FETCH_EXECUTE(0),TALU_OUTPUT,TALU_COUT);
--cont_alu_op,t_cin,
--talu_output,
--talu_cout); 

-- DecExc_input(24 DOWNTO 17),DecExc_input(16 DOWNTO 9),CONT_ALU_OP,T_CIN,tALU_OUTPUT,tALU_COUT);
WriteBack_Input<=talu_output&t_FETCH_EXECUTE(4 DOWNTO 2)&t_FETCH_EXECUTE(1);
--WriteBack register PORT MAP
-- writeback_mem: A_REGISTER GENERIC MAP (25) PORT MAP(tALU_OUTPUT,CLK,EN,RST,tWRITE_BACK_REGISTER);  
writeback_mem: A_REGISTER GENERIC MAP (12) PORT MAP(WriteBack_Input,CLK,EN,RST,tWRITE_BACK_REGISTER);  
tWRITE_PORT<=tWRITE_BACK_REGISTER(11 DOWNTO 4);
--WRITEBACK_ENABLE<=WriteBack_Input(0);
WRITEBACK_ENABLE<=tWRITE_BACK_REGISTER(0);
tWRITEBACK_ADDRESS<=tWRITE_BACK_REGISTER(3 DOWNTO 1);

--for the tWRITEBACK_ADDRESS signal we will need a multiplexer to supply this input. It selects from either writeback_mem Register (signal tWRITE_BACK_REGISTER
--directly from the instruction cache (signal T_FETCH)

END ARC;
