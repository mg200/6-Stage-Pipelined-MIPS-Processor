
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY IF_ID IS 
PORT(
INSTRUCTION: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
INSTRUCTIONPLUSONE: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
i_PC: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
CLK,EN,RST: IN STD_LOGIC;
FLUSH: IN STD_LOGIC;
INSTUCTION_OUTPUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
if_idplus: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
IF_ID_PC: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END ENTITY;


ARCHITECTURE ARC OF IF_ID IS 
BEGIN
--SYNCHRONOUS BUFFER
PROCESS (CLK)
BEGIN
IF RISING_EDGE(CLK) AND EN='1' THEN 
IF RST='1' THEN 
INSTUCTION_OUTPUT<=(OTHERS=>'0');
if_idplus<=(OTHERS=>'0');
IF_ID_PC<=(OTHERS=>'0');
ELSE
INSTUCTION_OUTPUT<=INSTRUCTION;
if_idplus<=INSTRUCTIONPLUSONE;
IF_ID_PC<=i_PC;
END IF;
-- --ADDED ON 17/6/2023 FROM 35 TO 38 VERY suspicious
-- ELSIF RISING_EDGE(CLK) AND EN='0' AND FLUSH='1' THEN 
-- INSTUCTION_OUTPUT<=(OTHERS=>'0');
-- if_idplus<=(OTHERS=>'0');
-- IF_ID_PC<=(OTHERS=>'0');
END IF;
END PROCESS;

END ARC;