
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DcacheDataSelector IS 

PORT
(
    OPCODE:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    IF_ID_MOST_SIG: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    INTERRUPT: IN STD_LOGIC;
    CCR_REG_VALUES: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    PC: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    Piped_EXMEM_PC: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    NormalData: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    DataToCommit: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    -- ALuOutputorSP: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);

END ENTITY;



ARCHITECTURE ARC OF DcacheDataSelector IS 
BEGIN 
-- push call interrupt  in order
-- DataToCommit<=STD_LOGIC_VECTOR(TO_UNSIGNED(TO_INTEGER(UNSIGNED(PC))+1,DataToCommit'LENGTH)) WHEN  OPCODE="01100" ELSE 
DataToCommit<=STD_LOGIC_VECTOR(TO_UNSIGNED(TO_INTEGER(UNSIGNED(Piped_EXMEM_PC))+1,DataToCommit'LENGTH)) WHEN  OPCODE="01100" ELSE 
CCR_REG_VALUES&"000"&STD_LOGIC_VECTOR(TO_UNSIGNED(TO_INTEGER(UNSIGNED(PC(9 DOWNTO 0)))+1,10))  
WHEN (INTERRUPT='1' AND (IF_ID_MOST_SIG="00111" OR IF_ID_MOST_SIG="10010"))  ELSE --LDM and IADD
CCR_REG_VALUES&"000"&PC(9 DOWNTO 0) WHEN INTERRUPT='1' ELSE
NormalData;
END ARC;