Library ieee;
Use ieee.std_logic_1164.all;
USE IEEE.numeric_std.all;
use IEEE.math_real.all;
--USE WORK.mytrialpackage.all;

ENTITY PC IS
GENERIC(N: INTEGER:=8);
PORT(CLK: IN STD_LOGIC:='1';
COUNT: inOUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
EN: IN STD_LOGIC:='1';
RST: IN STD_LOGIC:='0'
);
END ENTITY;

ARCHITECTURE ARC OF PC IS 

BEGIN


PROCESS(CLK)
VARIABLE TEMP:INTEGER:=0;
VARIABLE ALL_ONES:STD_LOGIC_VECTOR(N-1 DOWNTO 0):=(OTHERS=>'1');
BEGIN
IF RISING_EDGE(CLK) THEN
IF rst='1' then
temp:=0 ;
elsif
EN='1' and rst='0' THEN
IF COUNT /=ALL_ONES THEN
TEMP:=TEMP+1;
ELSE --EN='1' AND COUNT=ALL_ONES THEN
TEMP:=0;
END IF;
END IF;
END IF;
COUNT<=STD_LOGIC_VECTOR(TO_UNSIGNED(TEMP,COUNT'LENGTH));
END PROCESS;

END ARC;
