Library ieee;
Use ieee.std_logic_1164.all;

ENTITY MEM_WB IS ---the name might be misleading as this is ONLY A BUFFER and NOT cache data memory
PORT(
CLK,EN,RST: IN STD_LOGIC;
INPUT_DATA:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
WRITE_EN: IN STD_LOGIC;
WRITE_ADDRESS: IN STD_LOGIC_VECTOR(2 DOWNTO 0);--the destination in the register file that has propagated through the ALU
WRITEBACK_DATA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);

END MEM_WB;


ARCHITECTURE ARC OF MEM_WB IS
COMPONENT A_REGISTER IS
GENERIC(N: INTEGER:=16);
PORT( 
D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
CLK,EN,RST: IN STD_LOGIC;
Q: OUT  STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;


--
SIGNAL tREGISTER_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN 

dataregister: A_Register GENERIC MAP(8) PORT MAP(INPUT_DATA,CLK,EN,RST,tREGISTER_DATA);

PROCESS (CLK)
BEGIN


END PROCESS;
END ARC; 


