
Library ieee;
Use ieee.std_logic_1164.all;

ENTITY ABUFFER IS
GENERIC (N: INTEGER:=3);
PORT(
DATA: IN STD_lOGIC_VECTOR((2**N)-1 DOWNTO 0);
CLK,EN,RST:IN STD_LOGIC;
Address_In: INOUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
CONTROL1: INOUT STD_LOGIC;
CONTROL2: INOUT STD_LOGIC;
OUTPUT: OUT STD_lOGIC_VECTOR((2**N)-1 DOWNTO 0)
--Address_OUT: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
);

END ENTITY;

ARCHITECTURE ARC OF ABUFFER IS
COMPONENT A_REGISTER IS
GENERIC(N: INTEGER:=16);
PORT( 
D: IN STd_LOGIC_VECTOR(N-1 DOWNTO 0);--input
CLK,EN,RST: IN STD_LOGIC;
Q: OUT  STd_LOGIC_VECTOR(N-1 DOWNTO 0));--output
END COMPONENT;
BEGIN

REGISTERMAP: A_REGISTER GENERIC MAP (8) PORT MAP(DATA,CLK,EN,RST,OUTPUT); 
END ARC;