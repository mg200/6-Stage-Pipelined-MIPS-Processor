Library ieee;
Use ieee.std_logic_1164.all;
USE IEEE.numeric_std.all;
use IEEE.math_real.all;

ENTITY SIGNALDELAYBUFFER IS
PORT(
CLK: IN STD_LOGIC;
EN: IN STD_LOGIC;
RST: IN STD_LOGIC;
MEMTOREG: IN STD_LOGIC;
REGWRITE: IN STD_LOGIC;
WRITEADDRESS: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
R_type_ALUOUTPUT: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
AluOp_IN: IN STD_LOGIC_VECTOR(4 DOWNTO 0);--ADDED ON 17/6/2023
MEMTOREG_OP: OUT STD_LOGIC;
REGWRITE_OP: OUT STD_LOGIC;
WRITEADDRESS_OP: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
R_type_ALUOUTPUT_OP: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
ALUOP_op: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END ENTITY;
--0011001000111111

ARCHITECTURE ARC OF SIGNALDELAYBUFFER IS 

BEGIN 

PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) AND EN='1' THEN 
IF RST='1' THEN 
MEMTOREG_OP<='0';
REGWRITE_OP<='0';
WRITEADDRESS_OP<="000";
R_type_ALUOUTPUT_OP<=(OTHERS=>'0');
ALUOP_op<=(OTHERS=>'0');
ELSE 
MEMTOREG_OP<=MEMTOREG;
REGWRITE_OP<=REGWRITE;
WRITEADDRESS_OP<=WRITEADDRESS;
R_type_ALUOUTPUT_OP<=R_type_ALUOUTPUT;
ALUOP_op<=AluOp_IN;
END IF;
END IF;
END PROCESS;

END ARC;
