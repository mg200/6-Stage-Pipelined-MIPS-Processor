LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY PC_Reg IS 
PORT(CLK,EN,RST: IN STD_LOGIC;
PC_INPUT: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
PC_OUTPUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END PC_Reg;


ARCHITECTURE ARC OF PC_Reg IS 

BEGIN
PROCESS(CLK)
BEGIN
IF EN='1' THEN
IF RISING_EDGE(CLK) THEN
IF RST='1' THEN
PC_OUTPUT<=(OTHERS=>'0');
ELSE
PC_OUTPUT<=PC_INPUT;
END IF;
END IF;
END IF;
END PROCESS;
END ARC;


