Library ieee;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Forwarding IS 
PORT(
    	--EX/MEM WB SIGNAL and Address IN MEMORY STAGE 1
WB_EX_MEM: IN STD_LOGIC;
WB_Address_EX_MEM: IN STD_LOGIC_VECTOR (2 DOWNTO 0);

  	--MEM/MEM WB SIGNAL and Address IN MEMORY STAGE 2
WB_MEM_MEM: IN STD_LOGIC;
WB_Address_MEM_MEM: IN STD_LOGIC_VECTOR (2 DOWNTO 0);

	--MEM/WB WB SIGNAL and Address IN WRITE BACK STAGE
WB_MEM_WB: IN STD_LOGIC;
WB_Address_MEM_WB: IN STD_LOGIC_VECTOR (2 DOWNTO 0);

	-- Adresses of RS , RT IN DECODE STAGE
RS_Address: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
RT_Address: IN STD_LOGIC_VECTOR (2 DOWNTO 0);


	--Selecting Parameters of ALU by selection of Forwarding 2-bit selectors
--FIRST_ALU_INPUT_SELECTOR OR SECOND_ALU_INPUT_SELECTOR
			--  00 OUTPUT OF READ DATA  FROM ID/EX BUFFER
			-- 01 SELECTING OUTPUT OF ALU FROM EX/MEM BUFFER
			-- 10 SELECTING OUTPUT OF ALU FROM MEM/MEM BUFFER  
			-- 11 SELECTING OUTPUT OF ALU FROM MEM/WB BUFFER  
FIRST_ALU_INPUT_SELECTOR: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
SECOND_ALU_INPUT_SELECTOR: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
);
END ENTITY;


ARCHITECTURE FORWARD OF Forwarding IS


SIGNAL RS_EX_MEM:  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL RS_MEM_MEM:  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL RS_MEM_WB:  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL RT_EX_MEM:  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL RT_MEM_MEM:  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL RT_MEM_WB:  STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN


FIRST_ALU_INPUT_SELECTOR <= "01" WHEN (WB_EX_MEM ='1') AND (WB_Address_EX_MEM = RS_Address)
			ELSE "10" WHEN (WB_MEM_MEM ='1') AND  (WB_Address_MEM_MEM = RS_Address)
			ELSE "11" WHEN (WB_MEM_WB = '1') AND (WB_Address_MEM_WB = RS_Address)
			ELSE "00";

SECOND_ALU_INPUT_SELECTOR <= "01" WHEN (WB_EX_MEM ='1') AND (WB_Address_EX_MEM = RT_Address)
			ELSE "10" WHEN (WB_MEM_MEM ='1') AND  (WB_Address_MEM_MEM = RT_Address)
			ELSE "11" WHEN (WB_MEM_WB = '1') AND (WB_Address_MEM_WB = RT_Address)
			ELSE "00";
	

END FORWARD;

