Library ieee;
Use ieee.std_logic_1164.all;
USE IEEE.numeric_std.all;
use IEEE.math_real.all;


--WORKING AND TESTED--

ENTITY DECODER_GENERIC IS
GENERIC(N:INTEGER:=5);--if we want a 3x8 decoder we give it 3 
PORT(
EN: IN STD_LOGIC;
INPUT: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
OUTPUT: OUT STD_LOGIC_VECTOR ((2**N)-1 DOWNTO 0)
);
END DECODER_GENERIC;

ARCHITECTURE ARC OF DECODER_GENERIC IS
BEGIN
PROCESS (INPUT,EN)
VARIABLE TEMP:STD_LOGIC_VECTOR((2**N)-1 DOWNTO 0);
BEGIN
TEMP:=(OTHERS=>'0');
IF EN='1' THEN
TEMP(TO_INTEGER(UNSIGNED(INPUT))):='1';--REMEMBER THAT A VARIABLE GETS AN IMMEDIATE VALUE
OUTPUT<=TEMP;
ELSE
OUTPUT<=TEMP;
END IF;
END PROCESS;
END ARC;



-- process(number)
-- begin
--     result <= (others => '0');
--     result(to_integer(unsigned(number))) <= '1';
-- end process;
--THIS IS THE WAY TO WRITE THE ABOVE CODE WITHOUT USING A VARIABLE--THIS MIGHT BE "MORE" SYNTHESIZABLE