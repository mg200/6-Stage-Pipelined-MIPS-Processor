Library ieee;
Use ieee.std_logic_1164.all;
USE IEEE.numeric_std.all;
use IEEE.math_real.all;
--USE WORK.mytrialpackage.all;



ENTITY RAM_GENERIC IS
GENERIC(
--ADD_WIDTH: INTEGER:=64;
ADD_WIDTH: INTEGER:=6;
 DATA_WIDTH:INTEGER:=8);
PORT(
DATA_IN: IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
-- ADDRESS: IN STD_LOGIC_VECTOR(log2_unsigned(ADD_WIDTH)-1 DOWNTO 0);
ADDRESS: IN STD_LOGIC_VECTOR(ADD_WIDTH-1 DOWNTO 0);
READ_WRITE: IN STD_LOGIC:='1';--DEFAULT IS 1 TO WRITE
CLK: IN STD_LOGIC;
DATAOUT: OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)
);
END RAM_GENERIC;




ARCHITECTURE ARC OF RAM_GENERIC IS 
--------COMPONENTS------
COMPONENT DECODER_GENERIC IS
GENERIC(N:INTEGER:=5);--if we want a 3x8 decoder we give it 3 
PORT(
EN: IN STD_LOGIC;
INPUT: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
OUTPUT: OUT STD_LOGIC_VECTOR ((2**N)-1 DOWNTO 0)
);
END COMPONENT;

-------END OF COMPONENTS-------
-- TYPE register_type IS ARRAY(0 TO 7) of STD_LOGIC_VECTOR (7 DOWNTO 0);
-- SIGNAL reg : register_type ;

-- TYPE RAM_TYPE IS ARRAY (0 TO ADD_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
TYPE RAM_TYPE IS ARRAY (0 TO (2**ADD_WIDTH)-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
SIGNAL RAM: RAM_TYPE:=(others=>(others=>'0'));--initialization of the RAM


-- --clock constant
-- constant clock_period:time:=100 ns;
-- SIGNAL TCLK: STD_LOGIC:='1';

---IT IS HERE THAT YOU DECLARE ALL SIGNALS, TYPES, COMPONENTS, CONSTANTS----
BEGIN --BEGINNING OF ARHCITECTURE
--PORT MAPS (IF ANY) ARE DONE HERE IN THIS AREA, OUTSIDE ANY PROCESS


-- tCLK<=NOT tCLK AFTER CLOCK_PERIOD/2;
-- PROCESS(Tclk)
-- BEGIN
-- tclk<=NOT tCLK AFTER CLOCK_PERIOD/2;
-- END PROCESS;
----the above process has any effect only if it is triggered in the process below it and tCLK is in the sensitivity list
--insteaf of CLK
--OTHER ARCHITECTURAL COMPONENTS


PROCESS (CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
    IF READ_WRITE='1' THEN
    RAM(TO_INTEGER(UNSIGNED(ADDRESS)))<=DATA_IN;
--END IF;
     ELSE 
    DATAOUT<=RAM(TO_INTEGER(UNSIGNED(ADDRESS)));
    END IF;
END IF;
END PROCESS;




END ARC;




--TO REMEMBER--
-- 1. A PROCESS IS A SEQUENTIAL BLOCK OF CODE THAT IS IMPLEMENTED CONCURRENTLY WITH THE REST OF THE 
-- BLOCKS BETWEEN BEGIN AND END OF THE ARCHITECTURE, INCLUDING WITH RESPECT TO OTHER BLOCKS
-- 2. 




