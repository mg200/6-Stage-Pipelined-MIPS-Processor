LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY CCR_Register IS 
PORT(CLK,EN,RST: IN STD_LOGIC;
CCR_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
CCR: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
);
END CCR_Register;

ARCHITECTURE ARC OF CCR_Register IS 


BEGIN
PROCESS(CLK,CCR_IN)
BEGIN
IF RST='1' THEN 
CCR<="000";
ELSE
-- ELSIF FALLING_EDGE(CLK) THEN
IF EN='1' THEN
CCR<=CCR_IN;
END IF;
END IF;
END PROCESS;
-- PROCESS(CLK)
-- BEGIN
-- IF RST='1' THEN 
-- CCR<="000";
-- ELSIF FALLING_EDGE(CLK) THEN
-- IF EN='1' THEN
-- CCR<=CCR_IN;
-- END IF;
-- END IF;
-- END PROCESS;
END ARC;
